--VHDL cheat sheet --

--Library and package declerations--
library IEEE;
