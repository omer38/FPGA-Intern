--VHDL cheat sheet --
